module top import pkg::*; #(
)(
);
endmodule
